module Adder(
    input [7:0] A, B,
    output [15:0] RESULT
);

assign RESULT = A + B;

endmodule
