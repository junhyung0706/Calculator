module testbench();

reg clk, reset;		    // 클럭과 리셋 신호 정의
reg [17:0] DIN;		    // 테스트할 데이터 입력
wire [15:0] RESULT;		// 계산기 모듈로부터의 결과값
wire NEG;		        // 계산 결과가 음수인지 나타내는 플래그

// Calculator 모듈 인스턴스화
Calculator Calculator_0(
    .clk(clk),
    .reset(reset),
    .DIN(DIN),
    .RESULT(RESULT),
    .NEG(NEG)
);

// 클럭 신호 생성: 매 5시간 단위마다 클럭 신호 반전
initial clk = 0;
always #5 clk = ~clk;

initial begin
    reset = 0;				                // 초기 리셋 상태는 0
    #10 reset = 1;				            // 10 시간 단위 후 리셋을 1로 설정
    #10 reset = 0;				            // 다시 리셋을 0으로 돌려 계산기 모듈이 작동하게 함
    DIN = 18'b00_00000000_00000000;		    // 첫 번째 테스트 데이터 (연산 코드 00: 덧셈, A=0, B=0)
    #10 DIN = 18'b00_00000000_01011101;	    // 두 번째 테스트 데이터 (연산 코드 00: 덧셈, A=0, B=93)
    #10 DIN = 18'b00_11000010_11110110;	    // 세 번째 테스트 데이터 (연산 코드 00: 덧셈, A=194, B=246)
    #10 DIN = 18'b01_11001100_00000000;	    // 네 번째 테스트 데이터 (연산 코드 01: 뺄셈, A=204, B=0)
    #10 DIN = 18'b10_10000110_01011001;	    // 다섯 번째 테스트 데이터 (연산 코드 10: 곱셈, A=134, B=89)
    #10 DIN = 18'b01_00110110_10011011;	    // 여섯 번째 테스트 데이터 (연산 코드 01: 뺄셈, A=54, B=155)
    #10 DIN = 18'b01_00010010_00000111;	    // 일곱 번째 테스트 데이터 (연산 코드 01: 뺄셈, A=18, B=7)
    #10 DIN = 18'b10_11010000_00000000;	    // 여덟 번째 테스트 데이터 (연산 코드 10: 곱셈, A=208, B=0)
    #10 DIN = 18'b00_01010101_10101010;	    // 아홉 번째 테스트 데이터 (연산 코드 00: 덧셈, A=85, B=170)
    #10 DIN = 18'b10_00000000_00000000;	    // 열 번째 테스트 데이터 (연산 코드 10: 곱셈, A=0, B=0)
    #10 DIN = 18'b00_00000000_00000000;	    // 마지막 테스트 데이터 (연산 코드 00: 덧셈, A=0, B=0, 연산을 재시작하기 위한 초기화)
    #200 $stop;				                // 충분한 시간이 지난 후 시뮬레이션 중지
end

endmodule
