module tb_alu();

reg clk, reset;
reg [7:0] A, B;                  		// 8비트 피연산자 A와 B
reg [1:0] OP_CODE;               	// 연산을 지정하는 2비트 연산 코드
wire [15:0] RESULT;              	// 연산 결과를 나타내는 16비트 출력
wire NEG;                        	// 연산 결과가 음수인 경우를 나타내는 플래그

// ALU 모듈 인스턴스화
ALU ALU_0(
    .A(A),
    .B(B),
    .OP_CODE(OP_CODE),
    .RESULT(RESULT),
    .NEG(NEG)
);

// 클럭 생성 로직
initial clk = 0;
always #5 clk = ~clk;            	// 매 5 단위 시간마다 클럭의 값을 반전

// 테스트 시퀀스
initial begin
    reset = 0;
    #10 reset = 1;              		// 초기에 리셋을 활성화
    #10 reset = 0;              		// 리셋을 해제
    
    // 연산 코드 00 (덧셈), A와 B 모두 0
    OP_CODE <= 2'b00;
    A <= 8'b00000000;
    B <= 8'b00000000;
    
    // 연산 코드 00 (덧셈), A = 0, B = 93
    #10
    OP_CODE <= 2'b00;
    A <= 8'b00000000;
    B <= 8'b01011101;
    
    // 연산 코드 00 (덧셈), A = 194, B = 246
    #10
    OP_CODE <= 2'b00;
    A <= 8'b11000010;
    B <= 8'b11110110;

    // 연산 코드 01 (뺄셈), A = 204, B = 0
    #10
    OP_CODE <= 2'b01;
    A <= 8'b11001100;
    B <= 8'b00000000;

    // 연산 코드 10 (곱셈), A = 134, B = 89
    #10
    OP_CODE <= 2'b10;
    A <= 8'b10000110;
    B <= 8'b01011001;

    // 연산 코드 01 (뺄셈), A = 54, B = 155
    #10
    OP_CODE <= 2'b01;
    A <= 8'b00110110;
    B <= 8'b10011011;
    
    // 연산 코드 10 (곱셈), A = 18, B = 7
    #10
    OP_CODE <= 2'b10;
    A <= 8'b00010010;
    B <= 8'b00000111;
    
    // 연산 코드 10 (곱셈), A = 208, B = 0
    #10
    OP_CODE <= 2'b10;
    A <= 8'b11010000;
    B <= 8'b00000000;
    
    // 연산 코드 00 (덧셈), A = 85, B = 170
    #10
    OP_CODE <= 2'b00;
    A <= 8'b01010101;
    B <= 8'b10101010;
    
    // 연산 코드 10 (곱셈), A와 B 모두 0
    #10
    OP_CODE <= 2'b10;
    A <= 8'b00000000;
    B <= 8'b00000000;
    
    // 연산 코드 00 (덧셈), A와 B 모두 0
    #10
    OP_CODE <= 2'b00;
    A <= 8'b00000000;
    B <= 8'b00000000;

    #200 $stop;                 // 시뮬레이션 정지
end

endmodule
